<sevenseg_decoder module extracted>