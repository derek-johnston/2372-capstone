<buzzer_one_shot module extracted>