<debounce_oneshot module extracted>