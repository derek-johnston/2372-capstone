<clk_en_div module extracted>