<display_mux2 module extracted>