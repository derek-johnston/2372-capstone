<shot_counter module extracted>