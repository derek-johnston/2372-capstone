<shot_fsm module extracted>